��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&#;K0���r�X�	�m��2�Fc\K���ث&d�f����){袋r����v��<��1���s���:"�ٔ��L5^Kz��&�Y��6��5��<�����z)+ه��:�a���o��з�/.�hD�A�z<�����	^�u�S�m��*1�T�j�F +���1ab3�X�DK=��:*}��Cکퟪ�xK�`�o�6{J�d*����ba��ݬM��4H-i��M�X���e���P¬bG��f�U#%ƣ�P-��":4փ�F�ڂ����  ��wP&�hN� j���@����ג�ҩN�a��^}�X�,1�qSr�T��.��4q�v��-"����Lڭ��o�a�����7vY�����\;^�fӭ=����h��r�`��jN�u\
�Z��i<}߮r�2�|f�$�ՄL�ъ�$Wdi��O~~�R�xȠD�Qg:�>�����V�	oS�b �n/1x�w�M+;ʹ��)Ff���<)6�4`E�/#~e(��8�5x8�c�^?N��D��Ϭ�T`���o�Չ���X!�#����t��ۄnF��,�����[��}�<��m�{ā�I�n�u"�UW��1���`U�ࠔP���RA��	/����8�O(�	��tE�Z�*.�@��I�pYG�s�T����t��c��]��j��Fg�����Q��LM
F���yڱ�Ƿ#��F��yG��z5s-��E�Ǥ�"�%��}L���N�� ����`O(0��Bp>	^��3"#�,�哿a�1FO�_�CZx��	'�)�o��������ߪ��puaO<�+��t�tq���p˼̓S؍V��MD�V���X��V{�������4�a��'Q�Lr��2�r`{�J �����H{�s,�5��g�z��_9;Hѭ��a';5`2�d0�<E�ά�w�/�����ph�r�_W9��+"���[��s1x� ���4��Fa�%��Z|RN i�}B0����-m��v�3
���$&�R��=���Tht�p��N�t�_��~�~0s�؂�KVC�Q��@�:]����:��E�[�� (��ɯ�ֺP>�~�\��y%��oO�_���-*��̟�D���f�+x�P�~p���k�����Xm3�|�|�!�(�<�p��w���R	x}�?::Pcߍ��/R/�*_J���;���?����~�=�@�oR��`��L�
���y��+�xV`}[�K�9�l��hF���b9ՔE6��v�G�=�{�A�c��*t���)��}s��\���ZV���Aӎ�����#=����܊Iù���g�����7�vI/�{Y��v�|�V2j�=BG��}|�w�����^f}����Jqve:Rm��0�q �zy�;��cVv9C�'m�R����K+�� i���Q��6��W����!=:�&2�������]l�Byk��">4���Y�Z�$I@O4�v�n����*7ҍ �&=Xy=;��a#_��&��u�D�Fy����ҷ�$:W��s�^�r��1��o'�}c�|����/_ď���.{Z��Ni��n R� JXjC��ϦC�'lz۵������L� �9>�:農�5�N�����hF>p�$5�k�Atug���%�X�6�B���%��G2��A�$�������0�2_� J>�טI�[��'5-��-��\~�+�zg� @��ݼ|�~��.�a^z97A�gD;���8�l���5H�m����p�����V�}�G�U�kk�(y ����"`��O��a���Ͳ�z��;W�gl��Cz������3_�kd!X�@k���~s�3�v�*/o��љ���p4G������*C��P~(��4��>�xJ@6_7ag	-���3�'�Tޙ���V�Ԭ��t7�R���h{O�b�
1y���=|Ka�w���+T�U���l���>=%���{��)�P���&ê��W�_Dxz��eЅ҈;_�K�xP����[��tt��3s�z��!�C۾1������)���2P<�������7\P�^�سA46��<8��C�~̙C�_0��%z���D�������Ku;pm�]��b&Jcinkn��\K'@H��1�}mð�RA�}�Wt��2g�#�W	��N�#
��d`�c���$��t���#Z��;�ԁ"A��~��>J����"�i�%!���'�K���Q����U�8=�]
&I ]y�*V��u@��LfN���2;��Sɧi/���ѷ���*Ũ5ώu��=+��5Q^o5�����z0:������Xb�P��l�kcx9s��Joy9*���K7]�����W(�"�j��{X�R�H�?�y�Z0u�p����&�r��B�d�)�4w#����o��f��옿�b#Oǎ�w�
�"�3��(
�栰f��U�/��E)�L}3�6L�iML:��D#�}��)�+��a�~j���k����2ǎ<�G�A��F���
L�3"M?� ��D�1$y�8Ϫ���7"�҉�����"@4\��]Չ�6���ܟfT�oV5�z���z��`!�	���ɤ��v�¢���,-I	ƅ�^8�<	��_������
��E�]?��@k���>�0�����Qbվ�B���:�|���3N|g�����*�b#�Ζ�Z�,JdK��{m��P��,O�2�R�C�F|q´�8�!�6�&c�:	J�g�2�ڞ��4	���~����>a�4PkK6��u��k�q�TK*��X|�%R�'W��e!�n��yr�+��|�o.1I'�9oto1x�*8X?)=��[��~!�li��D̪�A�`�~��P�����{�ǻ�Y�
�> or��(��1����^z�.*�8x	��$q.j��/l�*�^dv�ָ^Q
leE�-r��O�b��;G��"O��ZA���g>X6qT01���7j�L��.��ѻ�<��v����.%Q�ֽ���ɜpH����(�a�)���kN�Y�{6K�D����u�򁳊����P���h�����1'�ʪ?}��m�/0��=(�v	J���@ 
���wbn�w%c�b���`�"?���M�A�7-�~J�L�ё"N��M�5g�WH{ҵ1�s��$���[0H���ڋ����7 9�̅�֌���o�8���ֆ6/�	T+u��_u|s>���JGMJ6�㕢�A���J&"$#{m��%:����g�'�0S�j�/��_6Sd��gN�3�zq3k,�K��b�gd��b��\�(=�����g�Sz��}�b:��M�o����+����7�;��c�<Q4�$F�ބ�S`
Ei�e�ɘ�ƞ�'-?l�@����'V{*���b�^��4�E�EB���5r5����U�����ޥ�� ��e�#��Ԥ��,@0�(��gx^��������{ �{4V�@��ږ�'��M���9?� �L��W�{5������Z�ʙ��J_��wB(	k�ğ�1sg�ޢ?�]��6�P����N�i;H�'��v��\��<,��������k?��Mp06����琗{s�OГ�v=E;4��]�ьՕ��>�P&��ga��Ti���Q"��)f��Ɵq�s�^�荺AM>�w1�Xa�B� �I���s���.]٩[�wۚ�tfR	[��&6�Y)Q���~�����b�a����BA����#P�����9KM��6��
d�`�W�G��KTS������>Iy]b��Q4���uk7�]�H�{��P���u�\!<ڽi�8T>{��Hj�X����$�:.��c��1g���jG}�������t���֋�@`�H��057�x!.$~Ɇ���i�u�t�oa�C��L�J�$oKߟA�m|��p��NcR&�U�D&�B��ݥ�d?�U���� ��a��3c�r�n4��x�y���ԇ�J0+�M�f���+�NR��e��������dOCpʥ~ ����u�����4����+]��Q�]�J���O<�y�nA�T8NA���@��	��kǲ�g�xGm�����4�]-�yy=k�9�'�wd�&^�V�lQ�Qy��w����=h�&n�^b�y]:ll�ݝ&nʯ;��`�;�t��E��E�2lr���[�Y�ǛM;>����&Q���Ry?iz5*����NSOZא�ő2�ʻw�|a�n�(L�:��̾�D�T9!g���g>UG�9��^ؓ:�&��W_�.F%ۖ��H�^*�=���>�yT�#�9&"�<M�j�X��oݒ@��;���|���{��ɘShN�3�"��e/�Tu��SL��7����6IG��>�І��C�g���_l��KH�s|`��e��Eb0	n*���ѯpr~9���#���)�����bB���ў��"��)~����z@(u�C�z�!��]8p���G��/	�Q>b^�̦1�1=>��W����G��Bkg��\���b��1�8��9�W����)"�.ۨ�Ek/��*���=e͚�/R��mL�S�\a1ix�v��	����8���2��(%��	�Dr�,c7a0雄20ۨ{:0D��ߥ�����l�K��;��/��կ�R�z�&��*����'�s 4~�x�OK����GЪT�6��&�n�T�3ۅ0x�����!l��*������AMW