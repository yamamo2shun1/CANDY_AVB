// candy_avb_test_qsys.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module candy_avb_test_qsys (
		input  wire        clk_clk,                           //                         clk.clk
		output wire        codec_clk_clk,                     //                   codec_clk.clk
		input  wire [3:0]  eth_mii_rx_d,                      //                         eth.mii_rx_d
		input  wire        eth_mii_rx_dv,                     //                            .mii_rx_dv
		input  wire        eth_mii_rx_err,                    //                            .mii_rx_err
		output wire [3:0]  eth_mii_tx_d,                      //                            .mii_tx_d
		output wire        eth_mii_tx_en,                     //                            .mii_tx_en
		output wire        eth_mii_tx_err,                    //                            .mii_tx_err
		input  wire        eth_mii_crs,                       //                            .mii_crs
		input  wire        eth_mii_col,                       //                            .mii_col
		output wire        eth_clk_clk,                       //                     eth_clk.clk
		inout  wire        eth_interrupt_export,              //               eth_interrupt.export
		output wire        eth_mdio_mdc,                      //                    eth_mdio.mdc
		input  wire        eth_mdio_mdio_in,                  //                            .mdio_in
		output wire        eth_mdio_mdio_out,                 //                            .mdio_out
		output wire        eth_mdio_mdio_oen,                 //                            .mdio_oen
		input  wire        eth_misc_ff_tx_crc_fwd,            //                    eth_misc.ff_tx_crc_fwd
		output wire        eth_misc_ff_tx_septy,              //                            .ff_tx_septy
		output wire        eth_misc_tx_ff_uflow,              //                            .tx_ff_uflow
		output wire        eth_misc_ff_tx_a_full,             //                            .ff_tx_a_full
		output wire        eth_misc_ff_tx_a_empty,            //                            .ff_tx_a_empty
		output wire [17:0] eth_misc_rx_err_stat,              //                            .rx_err_stat
		output wire [3:0]  eth_misc_rx_frm_type,              //                            .rx_frm_type
		output wire        eth_misc_ff_rx_dsav,               //                            .ff_rx_dsav
		output wire        eth_misc_ff_rx_a_full,             //                            .ff_rx_a_full
		output wire        eth_misc_ff_rx_a_empty,            //                            .ff_rx_a_empty
		input  wire        eth_rx_clk_clk,                    //                  eth_rx_clk.clk
		input  wire        eth_status_set_10,                 //                  eth_status.set_10
		input  wire        eth_status_set_1000,               //                            .set_1000
		output wire        eth_status_eth_mode,               //                            .eth_mode
		output wire        eth_status_ena_10,                 //                            .ena_10
		input  wire        eth_tx_clk_clk,                    //                  eth_tx_clk.clk
		output wire [11:0] new_sdram_controller_0_wire_addr,  // new_sdram_controller_0_wire.addr
		output wire [1:0]  new_sdram_controller_0_wire_ba,    //                            .ba
		output wire        new_sdram_controller_0_wire_cas_n, //                            .cas_n
		output wire        new_sdram_controller_0_wire_cke,   //                            .cke
		output wire        new_sdram_controller_0_wire_cs_n,  //                            .cs_n
		inout  wire [15:0] new_sdram_controller_0_wire_dq,    //                            .dq
		output wire [1:0]  new_sdram_controller_0_wire_dqm,   //                            .dqm
		output wire        new_sdram_controller_0_wire_ras_n, //                            .ras_n
		output wire        new_sdram_controller_0_wire_we_n,  //                            .we_n
		input  wire        reset_reset_n,                     //                       reset.reset_n
		output wire        sdclk_clk_clk,                     //                   sdclk_clk.clk
		input  wire        uart0_rxd,                         //                       uart0.rxd
		output wire        uart0_txd,                         //                            .txd
		input  wire        uart0_cts_n,                       //                            .cts_n
		output wire        uart0_rts_n,                       //                            .rts_n
		output wire [1:0]  user_led_export                    //                    user_led.export
	);

	wire         tse_0_dma_tx_st_source_valid;                               // tse_0_dma_tx:st_source_valid -> tse_0_tse:ff_tx_wren
	wire  [31:0] tse_0_dma_tx_st_source_data;                                // tse_0_dma_tx:st_source_data -> tse_0_tse:ff_tx_data
	wire         tse_0_dma_tx_st_source_ready;                               // tse_0_tse:ff_tx_rdy -> tse_0_dma_tx:st_source_ready
	wire         tse_0_dma_tx_st_source_startofpacket;                       // tse_0_dma_tx:st_source_startofpacket -> tse_0_tse:ff_tx_sop
	wire         tse_0_dma_tx_st_source_endofpacket;                         // tse_0_dma_tx:st_source_endofpacket -> tse_0_tse:ff_tx_eop
	wire         tse_0_dma_tx_st_source_error;                               // tse_0_dma_tx:st_source_error -> tse_0_tse:ff_tx_err
	wire   [1:0] tse_0_dma_tx_st_source_empty;                               // tse_0_dma_tx:st_source_empty -> tse_0_tse:ff_tx_mod
	wire         altpll_0_c0_clk;                                            // altpll_0:c0 -> [descriptor_memory:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, jtaguart_0:clk, mm_interconnect_0:altpll_0_c0_clk, new_sdram_controller_0:clk, nios2_0:clk, onchip_flash_0:clock, pio_0:clk, pio_1:clk, rst_controller_001:clk, sysid_qsys_0:clock, timer_0:clk, timer_1:clk, timer_2:clk, tse_0_tse:clk, uart_0:clk]
	wire         altpll_0_c4_clk;                                            // altpll_0:c4 -> [avalon_st_adapter:in_clk_0_clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, mm_interconnect_0:altpll_0_c4_clk, rst_controller_002:clk, tse_0_dma_rx:clock_clk, tse_0_dma_tx:clock_clk, tse_0_tse:ff_rx_clk, tse_0_tse:ff_tx_clk]
	wire  [31:0] nios2_0_data_master_readdata;                               // mm_interconnect_0:nios2_0_data_master_readdata -> nios2_0:d_readdata
	wire         nios2_0_data_master_waitrequest;                            // mm_interconnect_0:nios2_0_data_master_waitrequest -> nios2_0:d_waitrequest
	wire         nios2_0_data_master_debugaccess;                            // nios2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_0_data_master_debugaccess
	wire  [24:0] nios2_0_data_master_address;                                // nios2_0:d_address -> mm_interconnect_0:nios2_0_data_master_address
	wire   [3:0] nios2_0_data_master_byteenable;                             // nios2_0:d_byteenable -> mm_interconnect_0:nios2_0_data_master_byteenable
	wire         nios2_0_data_master_read;                                   // nios2_0:d_read -> mm_interconnect_0:nios2_0_data_master_read
	wire         nios2_0_data_master_readdatavalid;                          // mm_interconnect_0:nios2_0_data_master_readdatavalid -> nios2_0:d_readdatavalid
	wire         nios2_0_data_master_write;                                  // nios2_0:d_write -> mm_interconnect_0:nios2_0_data_master_write
	wire  [31:0] nios2_0_data_master_writedata;                              // nios2_0:d_writedata -> mm_interconnect_0:nios2_0_data_master_writedata
	wire  [31:0] tse_0_dma_tx_descriptor_read_master_readdata;               // mm_interconnect_0:tse_0_dma_tx_descriptor_read_master_readdata -> tse_0_dma_tx:descriptor_read_master_readdata
	wire         tse_0_dma_tx_descriptor_read_master_waitrequest;            // mm_interconnect_0:tse_0_dma_tx_descriptor_read_master_waitrequest -> tse_0_dma_tx:descriptor_read_master_waitrequest
	wire  [24:0] tse_0_dma_tx_descriptor_read_master_address;                // tse_0_dma_tx:descriptor_read_master_address -> mm_interconnect_0:tse_0_dma_tx_descriptor_read_master_address
	wire         tse_0_dma_tx_descriptor_read_master_read;                   // tse_0_dma_tx:descriptor_read_master_read -> mm_interconnect_0:tse_0_dma_tx_descriptor_read_master_read
	wire         tse_0_dma_tx_descriptor_read_master_readdatavalid;          // mm_interconnect_0:tse_0_dma_tx_descriptor_read_master_readdatavalid -> tse_0_dma_tx:descriptor_read_master_readdatavalid
	wire   [3:0] tse_0_dma_tx_descriptor_read_master_burstcount;             // tse_0_dma_tx:descriptor_read_master_burstcount -> mm_interconnect_0:tse_0_dma_tx_descriptor_read_master_burstcount
	wire  [31:0] tse_0_dma_rx_descriptor_read_master_readdata;               // mm_interconnect_0:tse_0_dma_rx_descriptor_read_master_readdata -> tse_0_dma_rx:descriptor_read_master_readdata
	wire         tse_0_dma_rx_descriptor_read_master_waitrequest;            // mm_interconnect_0:tse_0_dma_rx_descriptor_read_master_waitrequest -> tse_0_dma_rx:descriptor_read_master_waitrequest
	wire  [24:0] tse_0_dma_rx_descriptor_read_master_address;                // tse_0_dma_rx:descriptor_read_master_address -> mm_interconnect_0:tse_0_dma_rx_descriptor_read_master_address
	wire         tse_0_dma_rx_descriptor_read_master_read;                   // tse_0_dma_rx:descriptor_read_master_read -> mm_interconnect_0:tse_0_dma_rx_descriptor_read_master_read
	wire         tse_0_dma_rx_descriptor_read_master_readdatavalid;          // mm_interconnect_0:tse_0_dma_rx_descriptor_read_master_readdatavalid -> tse_0_dma_rx:descriptor_read_master_readdatavalid
	wire   [3:0] tse_0_dma_rx_descriptor_read_master_burstcount;             // tse_0_dma_rx:descriptor_read_master_burstcount -> mm_interconnect_0:tse_0_dma_rx_descriptor_read_master_burstcount
	wire         tse_0_dma_tx_descriptor_write_master_waitrequest;           // mm_interconnect_0:tse_0_dma_tx_descriptor_write_master_waitrequest -> tse_0_dma_tx:descriptor_write_master_waitrequest
	wire  [24:0] tse_0_dma_tx_descriptor_write_master_address;               // tse_0_dma_tx:descriptor_write_master_address -> mm_interconnect_0:tse_0_dma_tx_descriptor_write_master_address
	wire   [3:0] tse_0_dma_tx_descriptor_write_master_byteenable;            // tse_0_dma_tx:descriptor_write_master_byteenable -> mm_interconnect_0:tse_0_dma_tx_descriptor_write_master_byteenable
	wire   [1:0] tse_0_dma_tx_descriptor_write_master_response;              // mm_interconnect_0:tse_0_dma_tx_descriptor_write_master_response -> tse_0_dma_tx:descriptor_write_master_response
	wire         tse_0_dma_tx_descriptor_write_master_write;                 // tse_0_dma_tx:descriptor_write_master_write -> mm_interconnect_0:tse_0_dma_tx_descriptor_write_master_write
	wire  [31:0] tse_0_dma_tx_descriptor_write_master_writedata;             // tse_0_dma_tx:descriptor_write_master_writedata -> mm_interconnect_0:tse_0_dma_tx_descriptor_write_master_writedata
	wire         tse_0_dma_tx_descriptor_write_master_writeresponsevalid;    // mm_interconnect_0:tse_0_dma_tx_descriptor_write_master_writeresponsevalid -> tse_0_dma_tx:descriptor_write_master_writeresponsevalid
	wire         tse_0_dma_rx_descriptor_write_master_waitrequest;           // mm_interconnect_0:tse_0_dma_rx_descriptor_write_master_waitrequest -> tse_0_dma_rx:descriptor_write_master_waitrequest
	wire  [24:0] tse_0_dma_rx_descriptor_write_master_address;               // tse_0_dma_rx:descriptor_write_master_address -> mm_interconnect_0:tse_0_dma_rx_descriptor_write_master_address
	wire   [3:0] tse_0_dma_rx_descriptor_write_master_byteenable;            // tse_0_dma_rx:descriptor_write_master_byteenable -> mm_interconnect_0:tse_0_dma_rx_descriptor_write_master_byteenable
	wire   [1:0] tse_0_dma_rx_descriptor_write_master_response;              // mm_interconnect_0:tse_0_dma_rx_descriptor_write_master_response -> tse_0_dma_rx:descriptor_write_master_response
	wire         tse_0_dma_rx_descriptor_write_master_write;                 // tse_0_dma_rx:descriptor_write_master_write -> mm_interconnect_0:tse_0_dma_rx_descriptor_write_master_write
	wire  [31:0] tse_0_dma_rx_descriptor_write_master_writedata;             // tse_0_dma_rx:descriptor_write_master_writedata -> mm_interconnect_0:tse_0_dma_rx_descriptor_write_master_writedata
	wire         tse_0_dma_rx_descriptor_write_master_writeresponsevalid;    // mm_interconnect_0:tse_0_dma_rx_descriptor_write_master_writeresponsevalid -> tse_0_dma_rx:descriptor_write_master_writeresponsevalid
	wire  [31:0] nios2_0_instruction_master_readdata;                        // mm_interconnect_0:nios2_0_instruction_master_readdata -> nios2_0:i_readdata
	wire         nios2_0_instruction_master_waitrequest;                     // mm_interconnect_0:nios2_0_instruction_master_waitrequest -> nios2_0:i_waitrequest
	wire  [24:0] nios2_0_instruction_master_address;                         // nios2_0:i_address -> mm_interconnect_0:nios2_0_instruction_master_address
	wire         nios2_0_instruction_master_read;                            // nios2_0:i_read -> mm_interconnect_0:nios2_0_instruction_master_read
	wire         nios2_0_instruction_master_readdatavalid;                   // mm_interconnect_0:nios2_0_instruction_master_readdatavalid -> nios2_0:i_readdatavalid
	wire  [31:0] tse_0_dma_tx_mm_read_readdata;                              // mm_interconnect_0:tse_0_dma_tx_mm_read_readdata -> tse_0_dma_tx:mm_read_readdata
	wire         tse_0_dma_tx_mm_read_waitrequest;                           // mm_interconnect_0:tse_0_dma_tx_mm_read_waitrequest -> tse_0_dma_tx:mm_read_waitrequest
	wire  [23:0] tse_0_dma_tx_mm_read_address;                               // tse_0_dma_tx:mm_read_address -> mm_interconnect_0:tse_0_dma_tx_mm_read_address
	wire         tse_0_dma_tx_mm_read_read;                                  // tse_0_dma_tx:mm_read_read -> mm_interconnect_0:tse_0_dma_tx_mm_read_read
	wire   [3:0] tse_0_dma_tx_mm_read_byteenable;                            // tse_0_dma_tx:mm_read_byteenable -> mm_interconnect_0:tse_0_dma_tx_mm_read_byteenable
	wire         tse_0_dma_tx_mm_read_readdatavalid;                         // mm_interconnect_0:tse_0_dma_tx_mm_read_readdatavalid -> tse_0_dma_tx:mm_read_readdatavalid
	wire   [5:0] tse_0_dma_tx_mm_read_burstcount;                            // tse_0_dma_tx:mm_read_burstcount -> mm_interconnect_0:tse_0_dma_tx_mm_read_burstcount
	wire         tse_0_dma_rx_mm_write_waitrequest;                          // mm_interconnect_0:tse_0_dma_rx_mm_write_waitrequest -> tse_0_dma_rx:mm_write_waitrequest
	wire  [23:0] tse_0_dma_rx_mm_write_address;                              // tse_0_dma_rx:mm_write_address -> mm_interconnect_0:tse_0_dma_rx_mm_write_address
	wire   [3:0] tse_0_dma_rx_mm_write_byteenable;                           // tse_0_dma_rx:mm_write_byteenable -> mm_interconnect_0:tse_0_dma_rx_mm_write_byteenable
	wire         tse_0_dma_rx_mm_write_write;                                // tse_0_dma_rx:mm_write_write -> mm_interconnect_0:tse_0_dma_rx_mm_write_write
	wire  [31:0] tse_0_dma_rx_mm_write_writedata;                            // tse_0_dma_rx:mm_write_writedata -> mm_interconnect_0:tse_0_dma_rx_mm_write_writedata
	wire   [5:0] tse_0_dma_rx_mm_write_burstcount;                           // tse_0_dma_rx:mm_write_burstcount -> mm_interconnect_0:tse_0_dma_rx_mm_write_burstcount
	wire         mm_interconnect_0_jtaguart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtaguart_0_avalon_jtag_slave_chipselect -> jtaguart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtaguart_0_avalon_jtag_slave_readdata;    // jtaguart_0:av_readdata -> mm_interconnect_0:jtaguart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtaguart_0_avalon_jtag_slave_waitrequest; // jtaguart_0:av_waitrequest -> mm_interconnect_0:jtaguart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtaguart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtaguart_0_avalon_jtag_slave_address -> jtaguart_0:av_address
	wire         mm_interconnect_0_jtaguart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtaguart_0_avalon_jtag_slave_read -> jtaguart_0:av_read_n
	wire         mm_interconnect_0_jtaguart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtaguart_0_avalon_jtag_slave_write -> jtaguart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtaguart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtaguart_0_avalon_jtag_slave_writedata -> jtaguart_0:av_writedata
	wire  [31:0] mm_interconnect_0_tse_0_tse_control_port_readdata;          // tse_0_tse:reg_data_out -> mm_interconnect_0:tse_0_tse_control_port_readdata
	wire         mm_interconnect_0_tse_0_tse_control_port_waitrequest;       // tse_0_tse:reg_busy -> mm_interconnect_0:tse_0_tse_control_port_waitrequest
	wire   [7:0] mm_interconnect_0_tse_0_tse_control_port_address;           // mm_interconnect_0:tse_0_tse_control_port_address -> tse_0_tse:reg_addr
	wire         mm_interconnect_0_tse_0_tse_control_port_read;              // mm_interconnect_0:tse_0_tse_control_port_read -> tse_0_tse:reg_rd
	wire         mm_interconnect_0_tse_0_tse_control_port_write;             // mm_interconnect_0:tse_0_tse_control_port_write -> tse_0_tse:reg_wr
	wire  [31:0] mm_interconnect_0_tse_0_tse_control_port_writedata;         // mm_interconnect_0:tse_0_tse_control_port_writedata -> tse_0_tse:reg_data_in
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;      // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;       // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_tse_0_dma_rx_csr_readdata;                // tse_0_dma_rx:csr_readdata -> mm_interconnect_0:tse_0_dma_rx_csr_readdata
	wire   [2:0] mm_interconnect_0_tse_0_dma_rx_csr_address;                 // mm_interconnect_0:tse_0_dma_rx_csr_address -> tse_0_dma_rx:csr_address
	wire         mm_interconnect_0_tse_0_dma_rx_csr_read;                    // mm_interconnect_0:tse_0_dma_rx_csr_read -> tse_0_dma_rx:csr_read
	wire   [3:0] mm_interconnect_0_tse_0_dma_rx_csr_byteenable;              // mm_interconnect_0:tse_0_dma_rx_csr_byteenable -> tse_0_dma_rx:csr_byteenable
	wire         mm_interconnect_0_tse_0_dma_rx_csr_write;                   // mm_interconnect_0:tse_0_dma_rx_csr_write -> tse_0_dma_rx:csr_write
	wire  [31:0] mm_interconnect_0_tse_0_dma_rx_csr_writedata;               // mm_interconnect_0:tse_0_dma_rx_csr_writedata -> tse_0_dma_rx:csr_writedata
	wire  [31:0] mm_interconnect_0_tse_0_dma_tx_csr_readdata;                // tse_0_dma_tx:csr_readdata -> mm_interconnect_0:tse_0_dma_tx_csr_readdata
	wire   [2:0] mm_interconnect_0_tse_0_dma_tx_csr_address;                 // mm_interconnect_0:tse_0_dma_tx_csr_address -> tse_0_dma_tx:csr_address
	wire         mm_interconnect_0_tse_0_dma_tx_csr_read;                    // mm_interconnect_0:tse_0_dma_tx_csr_read -> tse_0_dma_tx:csr_read
	wire   [3:0] mm_interconnect_0_tse_0_dma_tx_csr_byteenable;              // mm_interconnect_0:tse_0_dma_tx_csr_byteenable -> tse_0_dma_tx:csr_byteenable
	wire         mm_interconnect_0_tse_0_dma_tx_csr_write;                   // mm_interconnect_0:tse_0_dma_tx_csr_write -> tse_0_dma_tx:csr_write
	wire  [31:0] mm_interconnect_0_tse_0_dma_tx_csr_writedata;               // mm_interconnect_0:tse_0_dma_tx_csr_writedata -> tse_0_dma_tx:csr_writedata
	wire  [31:0] mm_interconnect_0_onchip_flash_0_csr_readdata;              // onchip_flash_0:avmm_csr_readdata -> mm_interconnect_0:onchip_flash_0_csr_readdata
	wire   [0:0] mm_interconnect_0_onchip_flash_0_csr_address;               // mm_interconnect_0:onchip_flash_0_csr_address -> onchip_flash_0:avmm_csr_addr
	wire         mm_interconnect_0_onchip_flash_0_csr_read;                  // mm_interconnect_0:onchip_flash_0_csr_read -> onchip_flash_0:avmm_csr_read
	wire         mm_interconnect_0_onchip_flash_0_csr_write;                 // mm_interconnect_0:onchip_flash_0_csr_write -> onchip_flash_0:avmm_csr_write
	wire  [31:0] mm_interconnect_0_onchip_flash_0_csr_writedata;             // mm_interconnect_0:onchip_flash_0_csr_writedata -> onchip_flash_0:avmm_csr_writedata
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_readdata;             // onchip_flash_0:avmm_data_readdata -> mm_interconnect_0:onchip_flash_0_data_readdata
	wire         mm_interconnect_0_onchip_flash_0_data_waitrequest;          // onchip_flash_0:avmm_data_waitrequest -> mm_interconnect_0:onchip_flash_0_data_waitrequest
	wire  [15:0] mm_interconnect_0_onchip_flash_0_data_address;              // mm_interconnect_0:onchip_flash_0_data_address -> onchip_flash_0:avmm_data_addr
	wire         mm_interconnect_0_onchip_flash_0_data_read;                 // mm_interconnect_0:onchip_flash_0_data_read -> onchip_flash_0:avmm_data_read
	wire         mm_interconnect_0_onchip_flash_0_data_readdatavalid;        // onchip_flash_0:avmm_data_readdatavalid -> mm_interconnect_0:onchip_flash_0_data_readdatavalid
	wire         mm_interconnect_0_onchip_flash_0_data_write;                // mm_interconnect_0:onchip_flash_0_data_write -> onchip_flash_0:avmm_data_write
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_writedata;            // mm_interconnect_0:onchip_flash_0_data_writedata -> onchip_flash_0:avmm_data_writedata
	wire   [2:0] mm_interconnect_0_onchip_flash_0_data_burstcount;           // mm_interconnect_0:onchip_flash_0_data_burstcount -> onchip_flash_0:avmm_data_burstcount
	wire  [31:0] mm_interconnect_0_nios2_0_debug_mem_slave_readdata;         // nios2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_0_debug_mem_slave_waitrequest;      // nios2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_0_debug_mem_slave_debugaccess;      // mm_interconnect_0:nios2_0_debug_mem_slave_debugaccess -> nios2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_0_debug_mem_slave_address;          // mm_interconnect_0:nios2_0_debug_mem_slave_address -> nios2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_0_debug_mem_slave_read;             // mm_interconnect_0:nios2_0_debug_mem_slave_read -> nios2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_0_debug_mem_slave_byteenable;       // mm_interconnect_0:nios2_0_debug_mem_slave_byteenable -> nios2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_0_debug_mem_slave_write;            // mm_interconnect_0:nios2_0_debug_mem_slave_write -> nios2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_0_debug_mem_slave_writedata;        // mm_interconnect_0:nios2_0_debug_mem_slave_writedata -> nios2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;              // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;               // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                  // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                 // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;             // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire  [31:0] mm_interconnect_0_tse_0_dma_rx_prefetcher_csr_readdata;     // tse_0_dma_rx:prefetcher_csr_readdata -> mm_interconnect_0:tse_0_dma_rx_prefetcher_csr_readdata
	wire   [2:0] mm_interconnect_0_tse_0_dma_rx_prefetcher_csr_address;      // mm_interconnect_0:tse_0_dma_rx_prefetcher_csr_address -> tse_0_dma_rx:prefetcher_csr_address
	wire         mm_interconnect_0_tse_0_dma_rx_prefetcher_csr_read;         // mm_interconnect_0:tse_0_dma_rx_prefetcher_csr_read -> tse_0_dma_rx:prefetcher_csr_read
	wire         mm_interconnect_0_tse_0_dma_rx_prefetcher_csr_write;        // mm_interconnect_0:tse_0_dma_rx_prefetcher_csr_write -> tse_0_dma_rx:prefetcher_csr_write
	wire  [31:0] mm_interconnect_0_tse_0_dma_rx_prefetcher_csr_writedata;    // mm_interconnect_0:tse_0_dma_rx_prefetcher_csr_writedata -> tse_0_dma_rx:prefetcher_csr_writedata
	wire  [31:0] mm_interconnect_0_tse_0_dma_tx_prefetcher_csr_readdata;     // tse_0_dma_tx:prefetcher_csr_readdata -> mm_interconnect_0:tse_0_dma_tx_prefetcher_csr_readdata
	wire   [2:0] mm_interconnect_0_tse_0_dma_tx_prefetcher_csr_address;      // mm_interconnect_0:tse_0_dma_tx_prefetcher_csr_address -> tse_0_dma_tx:prefetcher_csr_address
	wire         mm_interconnect_0_tse_0_dma_tx_prefetcher_csr_read;         // mm_interconnect_0:tse_0_dma_tx_prefetcher_csr_read -> tse_0_dma_tx:prefetcher_csr_read
	wire         mm_interconnect_0_tse_0_dma_tx_prefetcher_csr_write;        // mm_interconnect_0:tse_0_dma_tx_prefetcher_csr_write -> tse_0_dma_tx:prefetcher_csr_write
	wire  [31:0] mm_interconnect_0_tse_0_dma_tx_prefetcher_csr_writedata;    // mm_interconnect_0:tse_0_dma_tx_prefetcher_csr_writedata -> tse_0_dma_tx:prefetcher_csr_writedata
	wire         mm_interconnect_0_pio_0_s1_chipselect;                      // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                        // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;                         // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;                           // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;                       // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire         mm_interconnect_0_uart_0_s1_chipselect;                     // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                       // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                        // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;                           // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                  // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;                          // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                      // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         mm_interconnect_0_timer_1_s1_chipselect;                    // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                      // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                       // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                         // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                     // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                    // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                      // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                       // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                         // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                     // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_timer_2_s1_chipselect;                    // mm_interconnect_0:timer_2_s1_chipselect -> timer_2:chipselect
	wire  [15:0] mm_interconnect_0_timer_2_s1_readdata;                      // timer_2:readdata -> mm_interconnect_0:timer_2_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_2_s1_address;                       // mm_interconnect_0:timer_2_s1_address -> timer_2:address
	wire         mm_interconnect_0_timer_2_s1_write;                         // mm_interconnect_0:timer_2_s1_write -> timer_2:write_n
	wire  [15:0] mm_interconnect_0_timer_2_s1_writedata;                     // mm_interconnect_0:timer_2_s1_writedata -> timer_2:writedata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_chipselect;     // mm_interconnect_0:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	wire  [15:0] mm_interconnect_0_new_sdram_controller_0_s1_readdata;       // new_sdram_controller_0:za_data -> mm_interconnect_0:new_sdram_controller_0_s1_readdata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_waitrequest;    // new_sdram_controller_0:za_waitrequest -> mm_interconnect_0:new_sdram_controller_0_s1_waitrequest
	wire  [21:0] mm_interconnect_0_new_sdram_controller_0_s1_address;        // mm_interconnect_0:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	wire         mm_interconnect_0_new_sdram_controller_0_s1_read;           // mm_interconnect_0:new_sdram_controller_0_s1_read -> new_sdram_controller_0:az_rd_n
	wire   [1:0] mm_interconnect_0_new_sdram_controller_0_s1_byteenable;     // mm_interconnect_0:new_sdram_controller_0_s1_byteenable -> new_sdram_controller_0:az_be_n
	wire         mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid;  // new_sdram_controller_0:za_valid -> mm_interconnect_0:new_sdram_controller_0_s1_readdatavalid
	wire         mm_interconnect_0_new_sdram_controller_0_s1_write;          // mm_interconnect_0:new_sdram_controller_0_s1_write -> new_sdram_controller_0:az_wr_n
	wire  [15:0] mm_interconnect_0_new_sdram_controller_0_s1_writedata;      // mm_interconnect_0:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	wire         mm_interconnect_0_pio_1_s1_chipselect;                      // mm_interconnect_0:pio_1_s1_chipselect -> pio_1:chipselect
	wire  [31:0] mm_interconnect_0_pio_1_s1_readdata;                        // pio_1:readdata -> mm_interconnect_0:pio_1_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_1_s1_address;                         // mm_interconnect_0:pio_1_s1_address -> pio_1:address
	wire         mm_interconnect_0_pio_1_s1_write;                           // mm_interconnect_0:pio_1_s1_write -> pio_1:write_n
	wire  [31:0] mm_interconnect_0_pio_1_s1_writedata;                       // mm_interconnect_0:pio_1_s1_writedata -> pio_1:writedata
	wire         mm_interconnect_0_descriptor_memory_s1_chipselect;          // mm_interconnect_0:descriptor_memory_s1_chipselect -> descriptor_memory:chipselect
	wire  [31:0] mm_interconnect_0_descriptor_memory_s1_readdata;            // descriptor_memory:readdata -> mm_interconnect_0:descriptor_memory_s1_readdata
	wire   [9:0] mm_interconnect_0_descriptor_memory_s1_address;             // mm_interconnect_0:descriptor_memory_s1_address -> descriptor_memory:address
	wire   [3:0] mm_interconnect_0_descriptor_memory_s1_byteenable;          // mm_interconnect_0:descriptor_memory_s1_byteenable -> descriptor_memory:byteenable
	wire         mm_interconnect_0_descriptor_memory_s1_write;               // mm_interconnect_0:descriptor_memory_s1_write -> descriptor_memory:write
	wire  [31:0] mm_interconnect_0_descriptor_memory_s1_writedata;           // mm_interconnect_0:descriptor_memory_s1_writedata -> descriptor_memory:writedata
	wire         mm_interconnect_0_descriptor_memory_s1_clken;               // mm_interconnect_0:descriptor_memory_s1_clken -> descriptor_memory:clken
	wire         irq_mapper_receiver2_irq;                                   // jtaguart_0:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                   // uart_0:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                   // timer_0:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                   // timer_1:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                   // timer_2:irq -> irq_mapper:receiver6_irq
	wire  [31:0] nios2_0_irq_irq;                                            // irq_mapper:sender_irq -> nios2_0:irq
	wire         irq_mapper_receiver0_irq;                                   // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                              // tse_0_dma_tx:csr_irq_irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                   // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                          // tse_0_dma_rx:csr_irq_irq -> irq_synchronizer_001:receiver_irq
	wire         tse_0_tse_receive_valid;                                    // tse_0_tse:ff_rx_dval -> avalon_st_adapter:in_0_valid
	wire  [31:0] tse_0_tse_receive_data;                                     // tse_0_tse:ff_rx_data -> avalon_st_adapter:in_0_data
	wire         tse_0_tse_receive_ready;                                    // avalon_st_adapter:in_0_ready -> tse_0_tse:ff_rx_rdy
	wire         tse_0_tse_receive_startofpacket;                            // tse_0_tse:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	wire         tse_0_tse_receive_endofpacket;                              // tse_0_tse:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	wire   [5:0] tse_0_tse_receive_error;                                    // tse_0_tse:rx_err -> avalon_st_adapter:in_0_error
	wire   [1:0] tse_0_tse_receive_empty;                                    // tse_0_tse:ff_rx_mod -> avalon_st_adapter:in_0_empty
	wire         avalon_st_adapter_out_0_valid;                              // avalon_st_adapter:out_0_valid -> tse_0_dma_rx:st_sink_valid
	wire  [31:0] avalon_st_adapter_out_0_data;                               // avalon_st_adapter:out_0_data -> tse_0_dma_rx:st_sink_data
	wire         avalon_st_adapter_out_0_ready;                              // tse_0_dma_rx:st_sink_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                      // avalon_st_adapter:out_0_startofpacket -> tse_0_dma_rx:st_sink_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                        // avalon_st_adapter:out_0_endofpacket -> tse_0_dma_rx:st_sink_endofpacket
	wire   [5:0] avalon_st_adapter_out_0_error;                              // avalon_st_adapter:out_0_error -> tse_0_dma_rx:st_sink_error
	wire   [1:0] avalon_st_adapter_out_0_empty;                              // avalon_st_adapter:out_0_empty -> tse_0_dma_rx:st_sink_empty
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         nios2_0_debug_reset_request_reset;                          // nios2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> [descriptor_memory:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, jtaguart_0:rst_n, mm_interconnect_0:nios2_0_reset_reset_bridge_in_reset_reset, new_sdram_controller_0:reset_n, nios2_0:reset_n, onchip_flash_0:reset_n, pio_0:reset_n, pio_1:reset_n, rst_translator:in_reset, sysid_qsys_0:reset_n, timer_0:reset_n, timer_1:reset_n, timer_2:reset_n, tse_0_tse:reset, uart_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                     // rst_controller_001:reset_req -> [descriptor_memory:reset_req, nios2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                         // rst_controller_002:reset_out -> [avalon_st_adapter:in_rst_0_reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, mm_interconnect_0:tse_0_dma_tx_reset_n_reset_bridge_in_reset_reset, tse_0_dma_rx:reset_n_reset_n, tse_0_dma_tx:reset_n_reset_n]

	candy_avb_test_qsys_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                 // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_0_c0_clk),                                //                    c0.clk
		.c1                 (sdclk_clk_clk),                                  //                    c1.clk
		.c2                 (codec_clk_clk),                                  //                    c2.clk
		.c3                 (eth_clk_clk),                                    //                    c3.clk
		.c4                 (altpll_0_c4_clk),                                //                    c4.clk
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.areset             (1'b0),                                           //           (terminated)
		.locked             (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (3'b000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	candy_avb_test_qsys_descriptor_memory descriptor_memory (
		.clk        (altpll_0_c0_clk),                                   //   clk1.clk
		.address    (mm_interconnect_0_descriptor_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_descriptor_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_descriptor_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_descriptor_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_descriptor_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_descriptor_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_descriptor_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                               // (terminated)
	);

	candy_avb_test_qsys_jtaguart_0 jtaguart_0 (
		.clk            (altpll_0_c0_clk),                                            //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                        //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtaguart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtaguart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtaguart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtaguart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtaguart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtaguart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtaguart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                    //               irq.irq
	);

	candy_avb_test_qsys_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (altpll_0_c0_clk),                                           //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                       // reset.reset_n
		.az_addr        (mm_interconnect_0_new_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_new_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_new_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_new_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_new_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_new_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (new_sdram_controller_0_wire_addr),                          //  wire.export
		.zs_ba          (new_sdram_controller_0_wire_ba),                            //      .export
		.zs_cas_n       (new_sdram_controller_0_wire_cas_n),                         //      .export
		.zs_cke         (new_sdram_controller_0_wire_cke),                           //      .export
		.zs_cs_n        (new_sdram_controller_0_wire_cs_n),                          //      .export
		.zs_dq          (new_sdram_controller_0_wire_dq),                            //      .export
		.zs_dqm         (new_sdram_controller_0_wire_dqm),                           //      .export
		.zs_ras_n       (new_sdram_controller_0_wire_ras_n),                         //      .export
		.zs_we_n        (new_sdram_controller_0_wire_we_n)                           //      .export
	);

	candy_avb_test_qsys_nios2_0 nios2_0 (
		.clk                                 (altpll_0_c0_clk),                                       //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                //                          .reset_req
		.d_address                           (nios2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                       // custom_instruction_master.readra
	);

	altera_onchip_flash #(
		.INIT_FILENAME                       (""),
		.INIT_FILENAME_SIM                   (""),
		.DEVICE_FAMILY                       ("MAX 10"),
		.PART_NAME                           ("10M16SAU169C8G"),
		.DEVICE_ID                           ("16"),
		.SECTOR1_START_ADDR                  (0),
		.SECTOR1_END_ADDR                    (4095),
		.SECTOR2_START_ADDR                  (4096),
		.SECTOR2_END_ADDR                    (8191),
		.SECTOR3_START_ADDR                  (8192),
		.SECTOR3_END_ADDR                    (47103),
		.SECTOR4_START_ADDR                  (0),
		.SECTOR4_END_ADDR                    (0),
		.SECTOR5_START_ADDR                  (0),
		.SECTOR5_END_ADDR                    (0),
		.MIN_VALID_ADDR                      (0),
		.MAX_VALID_ADDR                      (47103),
		.MIN_UFM_VALID_ADDR                  (0),
		.MAX_UFM_VALID_ADDR                  (47103),
		.SECTOR1_MAP                         (1),
		.SECTOR2_MAP                         (2),
		.SECTOR3_MAP                         (3),
		.SECTOR4_MAP                         (0),
		.SECTOR5_MAP                         (0),
		.ADDR_RANGE1_END_ADDR                (47103),
		.ADDR_RANGE2_END_ADDR                (47103),
		.ADDR_RANGE1_OFFSET                  (1024),
		.ADDR_RANGE2_OFFSET                  (0),
		.ADDR_RANGE3_OFFSET                  (0),
		.AVMM_DATA_ADDR_WIDTH                (16),
		.AVMM_DATA_DATA_WIDTH                (32),
		.AVMM_DATA_BURSTCOUNT_WIDTH          (3),
		.SECTOR_READ_PROTECTION_MODE         (24),
		.FLASH_SEQ_READ_DATA_COUNT           (4),
		.FLASH_ADDR_ALIGNMENT_BITS           (2),
		.FLASH_READ_CYCLE_MAX_INDEX          (4),
		.FLASH_RESET_CYCLE_MAX_INDEX         (25),
		.FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  (120),
		.FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX (35000000),
		.FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX (30500),
		.PARALLEL_MODE                       (1),
		.READ_AND_WRITE_MODE                 (1),
		.WRAPPING_BURST_MODE                 (0),
		.IS_DUAL_BOOT                        ("False"),
		.IS_ERAM_SKIP                        ("True"),
		.IS_COMPRESSED_IMAGE                 ("False")
	) onchip_flash_0 (
		.clock                   (altpll_0_c0_clk),                                     //    clk.clk
		.reset_n                 (~rst_controller_001_reset_out_reset),                 // nreset.reset_n
		.avmm_data_addr          (mm_interconnect_0_onchip_flash_0_data_address),       //   data.address
		.avmm_data_read          (mm_interconnect_0_onchip_flash_0_data_read),          //       .read
		.avmm_data_writedata     (mm_interconnect_0_onchip_flash_0_data_writedata),     //       .writedata
		.avmm_data_write         (mm_interconnect_0_onchip_flash_0_data_write),         //       .write
		.avmm_data_readdata      (mm_interconnect_0_onchip_flash_0_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (mm_interconnect_0_onchip_flash_0_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (mm_interconnect_0_onchip_flash_0_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (mm_interconnect_0_onchip_flash_0_data_burstcount),    //       .burstcount
		.avmm_csr_addr           (mm_interconnect_0_onchip_flash_0_csr_address),        //    csr.address
		.avmm_csr_read           (mm_interconnect_0_onchip_flash_0_csr_read),           //       .read
		.avmm_csr_writedata      (mm_interconnect_0_onchip_flash_0_csr_writedata),      //       .writedata
		.avmm_csr_write          (mm_interconnect_0_onchip_flash_0_csr_write),          //       .write
		.avmm_csr_readdata       (mm_interconnect_0_onchip_flash_0_csr_readdata)        //       .readdata
	);

	candy_avb_test_qsys_pio_0 pio_0 (
		.clk        (altpll_0_c0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.out_port   (user_led_export)                        // external_connection.export
	);

	candy_avb_test_qsys_pio_1 pio_1 (
		.clk        (altpll_0_c0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_0_pio_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_1_s1_readdata),   //                    .readdata
		.bidir_port (eth_interrupt_export)                   // external_connection.export
	);

	candy_avb_test_qsys_sysid_qsys_0 sysid_qsys_0 (
		.clock    (altpll_0_c0_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	candy_avb_test_qsys_timer_0 timer_0 (
		.clk        (altpll_0_c0_clk),                         //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)                 //   irq.irq
	);

	candy_avb_test_qsys_timer_0 timer_1 (
		.clk        (altpll_0_c0_clk),                         //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)                 //   irq.irq
	);

	candy_avb_test_qsys_timer_0 timer_2 (
		.clk        (altpll_0_c0_clk),                         //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_2_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_2_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_2_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_2_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_2_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver6_irq)                 //   irq.irq
	);

	candy_avb_test_qsys_tse_0_dma_rx tse_0_dma_rx (
		.mm_write_address                           (tse_0_dma_rx_mm_write_address),                           //                mm_write.address
		.mm_write_write                             (tse_0_dma_rx_mm_write_write),                             //                        .write
		.mm_write_byteenable                        (tse_0_dma_rx_mm_write_byteenable),                        //                        .byteenable
		.mm_write_writedata                         (tse_0_dma_rx_mm_write_writedata),                         //                        .writedata
		.mm_write_waitrequest                       (tse_0_dma_rx_mm_write_waitrequest),                       //                        .waitrequest
		.mm_write_burstcount                        (tse_0_dma_rx_mm_write_burstcount),                        //                        .burstcount
		.descriptor_read_master_address             (tse_0_dma_rx_descriptor_read_master_address),             //  descriptor_read_master.address
		.descriptor_read_master_read                (tse_0_dma_rx_descriptor_read_master_read),                //                        .read
		.descriptor_read_master_readdata            (tse_0_dma_rx_descriptor_read_master_readdata),            //                        .readdata
		.descriptor_read_master_waitrequest         (tse_0_dma_rx_descriptor_read_master_waitrequest),         //                        .waitrequest
		.descriptor_read_master_readdatavalid       (tse_0_dma_rx_descriptor_read_master_readdatavalid),       //                        .readdatavalid
		.descriptor_read_master_burstcount          (tse_0_dma_rx_descriptor_read_master_burstcount),          //                        .burstcount
		.descriptor_write_master_address            (tse_0_dma_rx_descriptor_write_master_address),            // descriptor_write_master.address
		.descriptor_write_master_write              (tse_0_dma_rx_descriptor_write_master_write),              //                        .write
		.descriptor_write_master_byteenable         (tse_0_dma_rx_descriptor_write_master_byteenable),         //                        .byteenable
		.descriptor_write_master_writedata          (tse_0_dma_rx_descriptor_write_master_writedata),          //                        .writedata
		.descriptor_write_master_waitrequest        (tse_0_dma_rx_descriptor_write_master_waitrequest),        //                        .waitrequest
		.descriptor_write_master_response           (tse_0_dma_rx_descriptor_write_master_response),           //                        .response
		.descriptor_write_master_writeresponsevalid (tse_0_dma_rx_descriptor_write_master_writeresponsevalid), //                        .writeresponsevalid
		.clock_clk                                  (altpll_0_c4_clk),                                         //                   clock.clk
		.reset_n_reset_n                            (~rst_controller_002_reset_out_reset),                     //                 reset_n.reset_n
		.csr_writedata                              (mm_interconnect_0_tse_0_dma_rx_csr_writedata),            //                     csr.writedata
		.csr_write                                  (mm_interconnect_0_tse_0_dma_rx_csr_write),                //                        .write
		.csr_byteenable                             (mm_interconnect_0_tse_0_dma_rx_csr_byteenable),           //                        .byteenable
		.csr_readdata                               (mm_interconnect_0_tse_0_dma_rx_csr_readdata),             //                        .readdata
		.csr_read                                   (mm_interconnect_0_tse_0_dma_rx_csr_read),                 //                        .read
		.csr_address                                (mm_interconnect_0_tse_0_dma_rx_csr_address),              //                        .address
		.prefetcher_csr_address                     (mm_interconnect_0_tse_0_dma_rx_prefetcher_csr_address),   //          prefetcher_csr.address
		.prefetcher_csr_read                        (mm_interconnect_0_tse_0_dma_rx_prefetcher_csr_read),      //                        .read
		.prefetcher_csr_write                       (mm_interconnect_0_tse_0_dma_rx_prefetcher_csr_write),     //                        .write
		.prefetcher_csr_writedata                   (mm_interconnect_0_tse_0_dma_rx_prefetcher_csr_writedata), //                        .writedata
		.prefetcher_csr_readdata                    (mm_interconnect_0_tse_0_dma_rx_prefetcher_csr_readdata),  //                        .readdata
		.csr_irq_irq                                (irq_synchronizer_001_receiver_irq),                       //                 csr_irq.irq
		.st_sink_data                               (avalon_st_adapter_out_0_data),                            //                 st_sink.data
		.st_sink_valid                              (avalon_st_adapter_out_0_valid),                           //                        .valid
		.st_sink_ready                              (avalon_st_adapter_out_0_ready),                           //                        .ready
		.st_sink_startofpacket                      (avalon_st_adapter_out_0_startofpacket),                   //                        .startofpacket
		.st_sink_endofpacket                        (avalon_st_adapter_out_0_endofpacket),                     //                        .endofpacket
		.st_sink_empty                              (avalon_st_adapter_out_0_empty),                           //                        .empty
		.st_sink_error                              (avalon_st_adapter_out_0_error)                            //                        .error
	);

	candy_avb_test_qsys_tse_0_dma_tx tse_0_dma_tx (
		.mm_read_address                            (tse_0_dma_tx_mm_read_address),                            //                 mm_read.address
		.mm_read_read                               (tse_0_dma_tx_mm_read_read),                               //                        .read
		.mm_read_byteenable                         (tse_0_dma_tx_mm_read_byteenable),                         //                        .byteenable
		.mm_read_readdata                           (tse_0_dma_tx_mm_read_readdata),                           //                        .readdata
		.mm_read_waitrequest                        (tse_0_dma_tx_mm_read_waitrequest),                        //                        .waitrequest
		.mm_read_readdatavalid                      (tse_0_dma_tx_mm_read_readdatavalid),                      //                        .readdatavalid
		.mm_read_burstcount                         (tse_0_dma_tx_mm_read_burstcount),                         //                        .burstcount
		.descriptor_read_master_address             (tse_0_dma_tx_descriptor_read_master_address),             //  descriptor_read_master.address
		.descriptor_read_master_read                (tse_0_dma_tx_descriptor_read_master_read),                //                        .read
		.descriptor_read_master_readdata            (tse_0_dma_tx_descriptor_read_master_readdata),            //                        .readdata
		.descriptor_read_master_waitrequest         (tse_0_dma_tx_descriptor_read_master_waitrequest),         //                        .waitrequest
		.descriptor_read_master_readdatavalid       (tse_0_dma_tx_descriptor_read_master_readdatavalid),       //                        .readdatavalid
		.descriptor_read_master_burstcount          (tse_0_dma_tx_descriptor_read_master_burstcount),          //                        .burstcount
		.descriptor_write_master_address            (tse_0_dma_tx_descriptor_write_master_address),            // descriptor_write_master.address
		.descriptor_write_master_write              (tse_0_dma_tx_descriptor_write_master_write),              //                        .write
		.descriptor_write_master_byteenable         (tse_0_dma_tx_descriptor_write_master_byteenable),         //                        .byteenable
		.descriptor_write_master_writedata          (tse_0_dma_tx_descriptor_write_master_writedata),          //                        .writedata
		.descriptor_write_master_waitrequest        (tse_0_dma_tx_descriptor_write_master_waitrequest),        //                        .waitrequest
		.descriptor_write_master_response           (tse_0_dma_tx_descriptor_write_master_response),           //                        .response
		.descriptor_write_master_writeresponsevalid (tse_0_dma_tx_descriptor_write_master_writeresponsevalid), //                        .writeresponsevalid
		.clock_clk                                  (altpll_0_c4_clk),                                         //                   clock.clk
		.reset_n_reset_n                            (~rst_controller_002_reset_out_reset),                     //                 reset_n.reset_n
		.csr_writedata                              (mm_interconnect_0_tse_0_dma_tx_csr_writedata),            //                     csr.writedata
		.csr_write                                  (mm_interconnect_0_tse_0_dma_tx_csr_write),                //                        .write
		.csr_byteenable                             (mm_interconnect_0_tse_0_dma_tx_csr_byteenable),           //                        .byteenable
		.csr_readdata                               (mm_interconnect_0_tse_0_dma_tx_csr_readdata),             //                        .readdata
		.csr_read                                   (mm_interconnect_0_tse_0_dma_tx_csr_read),                 //                        .read
		.csr_address                                (mm_interconnect_0_tse_0_dma_tx_csr_address),              //                        .address
		.prefetcher_csr_address                     (mm_interconnect_0_tse_0_dma_tx_prefetcher_csr_address),   //          prefetcher_csr.address
		.prefetcher_csr_read                        (mm_interconnect_0_tse_0_dma_tx_prefetcher_csr_read),      //                        .read
		.prefetcher_csr_write                       (mm_interconnect_0_tse_0_dma_tx_prefetcher_csr_write),     //                        .write
		.prefetcher_csr_writedata                   (mm_interconnect_0_tse_0_dma_tx_prefetcher_csr_writedata), //                        .writedata
		.prefetcher_csr_readdata                    (mm_interconnect_0_tse_0_dma_tx_prefetcher_csr_readdata),  //                        .readdata
		.csr_irq_irq                                (irq_synchronizer_receiver_irq),                           //                 csr_irq.irq
		.st_source_data                             (tse_0_dma_tx_st_source_data),                             //               st_source.data
		.st_source_valid                            (tse_0_dma_tx_st_source_valid),                            //                        .valid
		.st_source_ready                            (tse_0_dma_tx_st_source_ready),                            //                        .ready
		.st_source_startofpacket                    (tse_0_dma_tx_st_source_startofpacket),                    //                        .startofpacket
		.st_source_endofpacket                      (tse_0_dma_tx_st_source_endofpacket),                      //                        .endofpacket
		.st_source_empty                            (tse_0_dma_tx_st_source_empty),                            //                        .empty
		.st_source_error                            (tse_0_dma_tx_st_source_error)                             //                        .error
	);

	candy_avb_test_qsys_tse_0_tse tse_0_tse (
		.clk           (altpll_0_c0_clk),                                      // control_port_clock_connection.clk
		.reset         (rst_controller_001_reset_out_reset),                   //              reset_connection.reset
		.reg_addr      (mm_interconnect_0_tse_0_tse_control_port_address),     //                  control_port.address
		.reg_data_out  (mm_interconnect_0_tse_0_tse_control_port_readdata),    //                              .readdata
		.reg_rd        (mm_interconnect_0_tse_0_tse_control_port_read),        //                              .read
		.reg_data_in   (mm_interconnect_0_tse_0_tse_control_port_writedata),   //                              .writedata
		.reg_wr        (mm_interconnect_0_tse_0_tse_control_port_write),       //                              .write
		.reg_busy      (mm_interconnect_0_tse_0_tse_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (eth_tx_clk_clk),                                       //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (eth_rx_clk_clk),                                       //   pcs_mac_rx_clock_connection.clk
		.set_10        (eth_status_set_10),                                    //         mac_status_connection.set_10
		.set_1000      (eth_status_set_1000),                                  //                              .set_1000
		.eth_mode      (eth_status_eth_mode),                                  //                              .eth_mode
		.ena_10        (eth_status_ena_10),                                    //                              .ena_10
		.m_rx_d        (eth_mii_rx_d),                                         //            mac_mii_connection.mii_rx_d
		.m_rx_en       (eth_mii_rx_dv),                                        //                              .mii_rx_dv
		.m_rx_err      (eth_mii_rx_err),                                       //                              .mii_rx_err
		.m_tx_d        (eth_mii_tx_d),                                         //                              .mii_tx_d
		.m_tx_en       (eth_mii_tx_en),                                        //                              .mii_tx_en
		.m_tx_err      (eth_mii_tx_err),                                       //                              .mii_tx_err
		.m_rx_crs      (eth_mii_crs),                                          //                              .mii_crs
		.m_rx_col      (eth_mii_col),                                          //                              .mii_col
		.ff_rx_clk     (altpll_0_c4_clk),                                      //      receive_clock_connection.clk
		.ff_tx_clk     (altpll_0_c4_clk),                                      //     transmit_clock_connection.clk
		.ff_rx_data    (tse_0_tse_receive_data),                               //                       receive.data
		.ff_rx_eop     (tse_0_tse_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (tse_0_tse_receive_error),                              //                              .error
		.ff_rx_mod     (tse_0_tse_receive_empty),                              //                              .empty
		.ff_rx_rdy     (tse_0_tse_receive_ready),                              //                              .ready
		.ff_rx_sop     (tse_0_tse_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (tse_0_tse_receive_valid),                              //                              .valid
		.ff_tx_data    (tse_0_dma_tx_st_source_data),                          //                      transmit.data
		.ff_tx_eop     (tse_0_dma_tx_st_source_endofpacket),                   //                              .endofpacket
		.ff_tx_err     (tse_0_dma_tx_st_source_error),                         //                              .error
		.ff_tx_mod     (tse_0_dma_tx_st_source_empty),                         //                              .empty
		.ff_tx_rdy     (tse_0_dma_tx_st_source_ready),                         //                              .ready
		.ff_tx_sop     (tse_0_dma_tx_st_source_startofpacket),                 //                              .startofpacket
		.ff_tx_wren    (tse_0_dma_tx_st_source_valid),                         //                              .valid
		.mdc           (eth_mdio_mdc),                                         //           mac_mdio_connection.mdc
		.mdio_in       (eth_mdio_mdio_in),                                     //                              .mdio_in
		.mdio_out      (eth_mdio_mdio_out),                                    //                              .mdio_out
		.mdio_oen      (eth_mdio_mdio_oen),                                    //                              .mdio_oen
		.ff_tx_crc_fwd (eth_misc_ff_tx_crc_fwd),                               //           mac_misc_connection.ff_tx_crc_fwd
		.ff_tx_septy   (eth_misc_ff_tx_septy),                                 //                              .ff_tx_septy
		.tx_ff_uflow   (eth_misc_tx_ff_uflow),                                 //                              .tx_ff_uflow
		.ff_tx_a_full  (eth_misc_ff_tx_a_full),                                //                              .ff_tx_a_full
		.ff_tx_a_empty (eth_misc_ff_tx_a_empty),                               //                              .ff_tx_a_empty
		.rx_err_stat   (eth_misc_rx_err_stat),                                 //                              .rx_err_stat
		.rx_frm_type   (eth_misc_rx_frm_type),                                 //                              .rx_frm_type
		.ff_rx_dsav    (eth_misc_ff_rx_dsav),                                  //                              .ff_rx_dsav
		.ff_rx_a_full  (eth_misc_ff_rx_a_full),                                //                              .ff_rx_a_full
		.ff_rx_a_empty (eth_misc_ff_rx_a_empty)                                //                              .ff_rx_a_empty
	);

	candy_avb_test_qsys_uart_0 uart_0 (
		.clk           (altpll_0_c0_clk),                           //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.rxd           (uart0_rxd),                                 // external_connection.export
		.txd           (uart0_txd),                                 //                    .export
		.cts_n         (uart0_cts_n),                               //                    .export
		.rts_n         (uart0_rts_n),                               //                    .export
		.irq           (irq_mapper_receiver3_irq)                   //                 irq.irq
	);

	candy_avb_test_qsys_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                            (altpll_0_c0_clk),                                            //                                          altpll_0_c0.clk
		.altpll_0_c4_clk                                            (altpll_0_c4_clk),                                            //                                          altpll_0_c4.clk
		.clk_0_clk_clk                                              (clk_clk),                                                    //                                            clk_0_clk.clk
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2_0_reset_reset_bridge_in_reset_reset                  (rst_controller_001_reset_out_reset),                         //                  nios2_0_reset_reset_bridge_in_reset.reset
		.tse_0_dma_tx_reset_n_reset_bridge_in_reset_reset           (rst_controller_002_reset_out_reset),                         //           tse_0_dma_tx_reset_n_reset_bridge_in_reset.reset
		.nios2_0_data_master_address                                (nios2_0_data_master_address),                                //                                  nios2_0_data_master.address
		.nios2_0_data_master_waitrequest                            (nios2_0_data_master_waitrequest),                            //                                                     .waitrequest
		.nios2_0_data_master_byteenable                             (nios2_0_data_master_byteenable),                             //                                                     .byteenable
		.nios2_0_data_master_read                                   (nios2_0_data_master_read),                                   //                                                     .read
		.nios2_0_data_master_readdata                               (nios2_0_data_master_readdata),                               //                                                     .readdata
		.nios2_0_data_master_readdatavalid                          (nios2_0_data_master_readdatavalid),                          //                                                     .readdatavalid
		.nios2_0_data_master_write                                  (nios2_0_data_master_write),                                  //                                                     .write
		.nios2_0_data_master_writedata                              (nios2_0_data_master_writedata),                              //                                                     .writedata
		.nios2_0_data_master_debugaccess                            (nios2_0_data_master_debugaccess),                            //                                                     .debugaccess
		.nios2_0_instruction_master_address                         (nios2_0_instruction_master_address),                         //                           nios2_0_instruction_master.address
		.nios2_0_instruction_master_waitrequest                     (nios2_0_instruction_master_waitrequest),                     //                                                     .waitrequest
		.nios2_0_instruction_master_read                            (nios2_0_instruction_master_read),                            //                                                     .read
		.nios2_0_instruction_master_readdata                        (nios2_0_instruction_master_readdata),                        //                                                     .readdata
		.nios2_0_instruction_master_readdatavalid                   (nios2_0_instruction_master_readdatavalid),                   //                                                     .readdatavalid
		.tse_0_dma_rx_descriptor_read_master_address                (tse_0_dma_rx_descriptor_read_master_address),                //                  tse_0_dma_rx_descriptor_read_master.address
		.tse_0_dma_rx_descriptor_read_master_waitrequest            (tse_0_dma_rx_descriptor_read_master_waitrequest),            //                                                     .waitrequest
		.tse_0_dma_rx_descriptor_read_master_burstcount             (tse_0_dma_rx_descriptor_read_master_burstcount),             //                                                     .burstcount
		.tse_0_dma_rx_descriptor_read_master_read                   (tse_0_dma_rx_descriptor_read_master_read),                   //                                                     .read
		.tse_0_dma_rx_descriptor_read_master_readdata               (tse_0_dma_rx_descriptor_read_master_readdata),               //                                                     .readdata
		.tse_0_dma_rx_descriptor_read_master_readdatavalid          (tse_0_dma_rx_descriptor_read_master_readdatavalid),          //                                                     .readdatavalid
		.tse_0_dma_rx_descriptor_write_master_address               (tse_0_dma_rx_descriptor_write_master_address),               //                 tse_0_dma_rx_descriptor_write_master.address
		.tse_0_dma_rx_descriptor_write_master_waitrequest           (tse_0_dma_rx_descriptor_write_master_waitrequest),           //                                                     .waitrequest
		.tse_0_dma_rx_descriptor_write_master_byteenable            (tse_0_dma_rx_descriptor_write_master_byteenable),            //                                                     .byteenable
		.tse_0_dma_rx_descriptor_write_master_write                 (tse_0_dma_rx_descriptor_write_master_write),                 //                                                     .write
		.tse_0_dma_rx_descriptor_write_master_writedata             (tse_0_dma_rx_descriptor_write_master_writedata),             //                                                     .writedata
		.tse_0_dma_rx_descriptor_write_master_response              (tse_0_dma_rx_descriptor_write_master_response),              //                                                     .response
		.tse_0_dma_rx_descriptor_write_master_writeresponsevalid    (tse_0_dma_rx_descriptor_write_master_writeresponsevalid),    //                                                     .writeresponsevalid
		.tse_0_dma_rx_mm_write_address                              (tse_0_dma_rx_mm_write_address),                              //                                tse_0_dma_rx_mm_write.address
		.tse_0_dma_rx_mm_write_waitrequest                          (tse_0_dma_rx_mm_write_waitrequest),                          //                                                     .waitrequest
		.tse_0_dma_rx_mm_write_burstcount                           (tse_0_dma_rx_mm_write_burstcount),                           //                                                     .burstcount
		.tse_0_dma_rx_mm_write_byteenable                           (tse_0_dma_rx_mm_write_byteenable),                           //                                                     .byteenable
		.tse_0_dma_rx_mm_write_write                                (tse_0_dma_rx_mm_write_write),                                //                                                     .write
		.tse_0_dma_rx_mm_write_writedata                            (tse_0_dma_rx_mm_write_writedata),                            //                                                     .writedata
		.tse_0_dma_tx_descriptor_read_master_address                (tse_0_dma_tx_descriptor_read_master_address),                //                  tse_0_dma_tx_descriptor_read_master.address
		.tse_0_dma_tx_descriptor_read_master_waitrequest            (tse_0_dma_tx_descriptor_read_master_waitrequest),            //                                                     .waitrequest
		.tse_0_dma_tx_descriptor_read_master_burstcount             (tse_0_dma_tx_descriptor_read_master_burstcount),             //                                                     .burstcount
		.tse_0_dma_tx_descriptor_read_master_read                   (tse_0_dma_tx_descriptor_read_master_read),                   //                                                     .read
		.tse_0_dma_tx_descriptor_read_master_readdata               (tse_0_dma_tx_descriptor_read_master_readdata),               //                                                     .readdata
		.tse_0_dma_tx_descriptor_read_master_readdatavalid          (tse_0_dma_tx_descriptor_read_master_readdatavalid),          //                                                     .readdatavalid
		.tse_0_dma_tx_descriptor_write_master_address               (tse_0_dma_tx_descriptor_write_master_address),               //                 tse_0_dma_tx_descriptor_write_master.address
		.tse_0_dma_tx_descriptor_write_master_waitrequest           (tse_0_dma_tx_descriptor_write_master_waitrequest),           //                                                     .waitrequest
		.tse_0_dma_tx_descriptor_write_master_byteenable            (tse_0_dma_tx_descriptor_write_master_byteenable),            //                                                     .byteenable
		.tse_0_dma_tx_descriptor_write_master_write                 (tse_0_dma_tx_descriptor_write_master_write),                 //                                                     .write
		.tse_0_dma_tx_descriptor_write_master_writedata             (tse_0_dma_tx_descriptor_write_master_writedata),             //                                                     .writedata
		.tse_0_dma_tx_descriptor_write_master_response              (tse_0_dma_tx_descriptor_write_master_response),              //                                                     .response
		.tse_0_dma_tx_descriptor_write_master_writeresponsevalid    (tse_0_dma_tx_descriptor_write_master_writeresponsevalid),    //                                                     .writeresponsevalid
		.tse_0_dma_tx_mm_read_address                               (tse_0_dma_tx_mm_read_address),                               //                                 tse_0_dma_tx_mm_read.address
		.tse_0_dma_tx_mm_read_waitrequest                           (tse_0_dma_tx_mm_read_waitrequest),                           //                                                     .waitrequest
		.tse_0_dma_tx_mm_read_burstcount                            (tse_0_dma_tx_mm_read_burstcount),                            //                                                     .burstcount
		.tse_0_dma_tx_mm_read_byteenable                            (tse_0_dma_tx_mm_read_byteenable),                            //                                                     .byteenable
		.tse_0_dma_tx_mm_read_read                                  (tse_0_dma_tx_mm_read_read),                                  //                                                     .read
		.tse_0_dma_tx_mm_read_readdata                              (tse_0_dma_tx_mm_read_readdata),                              //                                                     .readdata
		.tse_0_dma_tx_mm_read_readdatavalid                         (tse_0_dma_tx_mm_read_readdatavalid),                         //                                                     .readdatavalid
		.altpll_0_pll_slave_address                                 (mm_interconnect_0_altpll_0_pll_slave_address),               //                                   altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                   (mm_interconnect_0_altpll_0_pll_slave_write),                 //                                                     .write
		.altpll_0_pll_slave_read                                    (mm_interconnect_0_altpll_0_pll_slave_read),                  //                                                     .read
		.altpll_0_pll_slave_readdata                                (mm_interconnect_0_altpll_0_pll_slave_readdata),              //                                                     .readdata
		.altpll_0_pll_slave_writedata                               (mm_interconnect_0_altpll_0_pll_slave_writedata),             //                                                     .writedata
		.descriptor_memory_s1_address                               (mm_interconnect_0_descriptor_memory_s1_address),             //                                 descriptor_memory_s1.address
		.descriptor_memory_s1_write                                 (mm_interconnect_0_descriptor_memory_s1_write),               //                                                     .write
		.descriptor_memory_s1_readdata                              (mm_interconnect_0_descriptor_memory_s1_readdata),            //                                                     .readdata
		.descriptor_memory_s1_writedata                             (mm_interconnect_0_descriptor_memory_s1_writedata),           //                                                     .writedata
		.descriptor_memory_s1_byteenable                            (mm_interconnect_0_descriptor_memory_s1_byteenable),          //                                                     .byteenable
		.descriptor_memory_s1_chipselect                            (mm_interconnect_0_descriptor_memory_s1_chipselect),          //                                                     .chipselect
		.descriptor_memory_s1_clken                                 (mm_interconnect_0_descriptor_memory_s1_clken),               //                                                     .clken
		.jtaguart_0_avalon_jtag_slave_address                       (mm_interconnect_0_jtaguart_0_avalon_jtag_slave_address),     //                         jtaguart_0_avalon_jtag_slave.address
		.jtaguart_0_avalon_jtag_slave_write                         (mm_interconnect_0_jtaguart_0_avalon_jtag_slave_write),       //                                                     .write
		.jtaguart_0_avalon_jtag_slave_read                          (mm_interconnect_0_jtaguart_0_avalon_jtag_slave_read),        //                                                     .read
		.jtaguart_0_avalon_jtag_slave_readdata                      (mm_interconnect_0_jtaguart_0_avalon_jtag_slave_readdata),    //                                                     .readdata
		.jtaguart_0_avalon_jtag_slave_writedata                     (mm_interconnect_0_jtaguart_0_avalon_jtag_slave_writedata),   //                                                     .writedata
		.jtaguart_0_avalon_jtag_slave_waitrequest                   (mm_interconnect_0_jtaguart_0_avalon_jtag_slave_waitrequest), //                                                     .waitrequest
		.jtaguart_0_avalon_jtag_slave_chipselect                    (mm_interconnect_0_jtaguart_0_avalon_jtag_slave_chipselect),  //                                                     .chipselect
		.new_sdram_controller_0_s1_address                          (mm_interconnect_0_new_sdram_controller_0_s1_address),        //                            new_sdram_controller_0_s1.address
		.new_sdram_controller_0_s1_write                            (mm_interconnect_0_new_sdram_controller_0_s1_write),          //                                                     .write
		.new_sdram_controller_0_s1_read                             (mm_interconnect_0_new_sdram_controller_0_s1_read),           //                                                     .read
		.new_sdram_controller_0_s1_readdata                         (mm_interconnect_0_new_sdram_controller_0_s1_readdata),       //                                                     .readdata
		.new_sdram_controller_0_s1_writedata                        (mm_interconnect_0_new_sdram_controller_0_s1_writedata),      //                                                     .writedata
		.new_sdram_controller_0_s1_byteenable                       (mm_interconnect_0_new_sdram_controller_0_s1_byteenable),     //                                                     .byteenable
		.new_sdram_controller_0_s1_readdatavalid                    (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid),  //                                                     .readdatavalid
		.new_sdram_controller_0_s1_waitrequest                      (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),    //                                                     .waitrequest
		.new_sdram_controller_0_s1_chipselect                       (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),     //                                                     .chipselect
		.nios2_0_debug_mem_slave_address                            (mm_interconnect_0_nios2_0_debug_mem_slave_address),          //                              nios2_0_debug_mem_slave.address
		.nios2_0_debug_mem_slave_write                              (mm_interconnect_0_nios2_0_debug_mem_slave_write),            //                                                     .write
		.nios2_0_debug_mem_slave_read                               (mm_interconnect_0_nios2_0_debug_mem_slave_read),             //                                                     .read
		.nios2_0_debug_mem_slave_readdata                           (mm_interconnect_0_nios2_0_debug_mem_slave_readdata),         //                                                     .readdata
		.nios2_0_debug_mem_slave_writedata                          (mm_interconnect_0_nios2_0_debug_mem_slave_writedata),        //                                                     .writedata
		.nios2_0_debug_mem_slave_byteenable                         (mm_interconnect_0_nios2_0_debug_mem_slave_byteenable),       //                                                     .byteenable
		.nios2_0_debug_mem_slave_waitrequest                        (mm_interconnect_0_nios2_0_debug_mem_slave_waitrequest),      //                                                     .waitrequest
		.nios2_0_debug_mem_slave_debugaccess                        (mm_interconnect_0_nios2_0_debug_mem_slave_debugaccess),      //                                                     .debugaccess
		.onchip_flash_0_csr_address                                 (mm_interconnect_0_onchip_flash_0_csr_address),               //                                   onchip_flash_0_csr.address
		.onchip_flash_0_csr_write                                   (mm_interconnect_0_onchip_flash_0_csr_write),                 //                                                     .write
		.onchip_flash_0_csr_read                                    (mm_interconnect_0_onchip_flash_0_csr_read),                  //                                                     .read
		.onchip_flash_0_csr_readdata                                (mm_interconnect_0_onchip_flash_0_csr_readdata),              //                                                     .readdata
		.onchip_flash_0_csr_writedata                               (mm_interconnect_0_onchip_flash_0_csr_writedata),             //                                                     .writedata
		.onchip_flash_0_data_address                                (mm_interconnect_0_onchip_flash_0_data_address),              //                                  onchip_flash_0_data.address
		.onchip_flash_0_data_write                                  (mm_interconnect_0_onchip_flash_0_data_write),                //                                                     .write
		.onchip_flash_0_data_read                                   (mm_interconnect_0_onchip_flash_0_data_read),                 //                                                     .read
		.onchip_flash_0_data_readdata                               (mm_interconnect_0_onchip_flash_0_data_readdata),             //                                                     .readdata
		.onchip_flash_0_data_writedata                              (mm_interconnect_0_onchip_flash_0_data_writedata),            //                                                     .writedata
		.onchip_flash_0_data_burstcount                             (mm_interconnect_0_onchip_flash_0_data_burstcount),           //                                                     .burstcount
		.onchip_flash_0_data_readdatavalid                          (mm_interconnect_0_onchip_flash_0_data_readdatavalid),        //                                                     .readdatavalid
		.onchip_flash_0_data_waitrequest                            (mm_interconnect_0_onchip_flash_0_data_waitrequest),          //                                                     .waitrequest
		.pio_0_s1_address                                           (mm_interconnect_0_pio_0_s1_address),                         //                                             pio_0_s1.address
		.pio_0_s1_write                                             (mm_interconnect_0_pio_0_s1_write),                           //                                                     .write
		.pio_0_s1_readdata                                          (mm_interconnect_0_pio_0_s1_readdata),                        //                                                     .readdata
		.pio_0_s1_writedata                                         (mm_interconnect_0_pio_0_s1_writedata),                       //                                                     .writedata
		.pio_0_s1_chipselect                                        (mm_interconnect_0_pio_0_s1_chipselect),                      //                                                     .chipselect
		.pio_1_s1_address                                           (mm_interconnect_0_pio_1_s1_address),                         //                                             pio_1_s1.address
		.pio_1_s1_write                                             (mm_interconnect_0_pio_1_s1_write),                           //                                                     .write
		.pio_1_s1_readdata                                          (mm_interconnect_0_pio_1_s1_readdata),                        //                                                     .readdata
		.pio_1_s1_writedata                                         (mm_interconnect_0_pio_1_s1_writedata),                       //                                                     .writedata
		.pio_1_s1_chipselect                                        (mm_interconnect_0_pio_1_s1_chipselect),                      //                                                     .chipselect
		.sysid_qsys_0_control_slave_address                         (mm_interconnect_0_sysid_qsys_0_control_slave_address),       //                           sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                        (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),      //                                                     .readdata
		.timer_0_s1_address                                         (mm_interconnect_0_timer_0_s1_address),                       //                                           timer_0_s1.address
		.timer_0_s1_write                                           (mm_interconnect_0_timer_0_s1_write),                         //                                                     .write
		.timer_0_s1_readdata                                        (mm_interconnect_0_timer_0_s1_readdata),                      //                                                     .readdata
		.timer_0_s1_writedata                                       (mm_interconnect_0_timer_0_s1_writedata),                     //                                                     .writedata
		.timer_0_s1_chipselect                                      (mm_interconnect_0_timer_0_s1_chipselect),                    //                                                     .chipselect
		.timer_1_s1_address                                         (mm_interconnect_0_timer_1_s1_address),                       //                                           timer_1_s1.address
		.timer_1_s1_write                                           (mm_interconnect_0_timer_1_s1_write),                         //                                                     .write
		.timer_1_s1_readdata                                        (mm_interconnect_0_timer_1_s1_readdata),                      //                                                     .readdata
		.timer_1_s1_writedata                                       (mm_interconnect_0_timer_1_s1_writedata),                     //                                                     .writedata
		.timer_1_s1_chipselect                                      (mm_interconnect_0_timer_1_s1_chipselect),                    //                                                     .chipselect
		.timer_2_s1_address                                         (mm_interconnect_0_timer_2_s1_address),                       //                                           timer_2_s1.address
		.timer_2_s1_write                                           (mm_interconnect_0_timer_2_s1_write),                         //                                                     .write
		.timer_2_s1_readdata                                        (mm_interconnect_0_timer_2_s1_readdata),                      //                                                     .readdata
		.timer_2_s1_writedata                                       (mm_interconnect_0_timer_2_s1_writedata),                     //                                                     .writedata
		.timer_2_s1_chipselect                                      (mm_interconnect_0_timer_2_s1_chipselect),                    //                                                     .chipselect
		.tse_0_dma_rx_csr_address                                   (mm_interconnect_0_tse_0_dma_rx_csr_address),                 //                                     tse_0_dma_rx_csr.address
		.tse_0_dma_rx_csr_write                                     (mm_interconnect_0_tse_0_dma_rx_csr_write),                   //                                                     .write
		.tse_0_dma_rx_csr_read                                      (mm_interconnect_0_tse_0_dma_rx_csr_read),                    //                                                     .read
		.tse_0_dma_rx_csr_readdata                                  (mm_interconnect_0_tse_0_dma_rx_csr_readdata),                //                                                     .readdata
		.tse_0_dma_rx_csr_writedata                                 (mm_interconnect_0_tse_0_dma_rx_csr_writedata),               //                                                     .writedata
		.tse_0_dma_rx_csr_byteenable                                (mm_interconnect_0_tse_0_dma_rx_csr_byteenable),              //                                                     .byteenable
		.tse_0_dma_rx_prefetcher_csr_address                        (mm_interconnect_0_tse_0_dma_rx_prefetcher_csr_address),      //                          tse_0_dma_rx_prefetcher_csr.address
		.tse_0_dma_rx_prefetcher_csr_write                          (mm_interconnect_0_tse_0_dma_rx_prefetcher_csr_write),        //                                                     .write
		.tse_0_dma_rx_prefetcher_csr_read                           (mm_interconnect_0_tse_0_dma_rx_prefetcher_csr_read),         //                                                     .read
		.tse_0_dma_rx_prefetcher_csr_readdata                       (mm_interconnect_0_tse_0_dma_rx_prefetcher_csr_readdata),     //                                                     .readdata
		.tse_0_dma_rx_prefetcher_csr_writedata                      (mm_interconnect_0_tse_0_dma_rx_prefetcher_csr_writedata),    //                                                     .writedata
		.tse_0_dma_tx_csr_address                                   (mm_interconnect_0_tse_0_dma_tx_csr_address),                 //                                     tse_0_dma_tx_csr.address
		.tse_0_dma_tx_csr_write                                     (mm_interconnect_0_tse_0_dma_tx_csr_write),                   //                                                     .write
		.tse_0_dma_tx_csr_read                                      (mm_interconnect_0_tse_0_dma_tx_csr_read),                    //                                                     .read
		.tse_0_dma_tx_csr_readdata                                  (mm_interconnect_0_tse_0_dma_tx_csr_readdata),                //                                                     .readdata
		.tse_0_dma_tx_csr_writedata                                 (mm_interconnect_0_tse_0_dma_tx_csr_writedata),               //                                                     .writedata
		.tse_0_dma_tx_csr_byteenable                                (mm_interconnect_0_tse_0_dma_tx_csr_byteenable),              //                                                     .byteenable
		.tse_0_dma_tx_prefetcher_csr_address                        (mm_interconnect_0_tse_0_dma_tx_prefetcher_csr_address),      //                          tse_0_dma_tx_prefetcher_csr.address
		.tse_0_dma_tx_prefetcher_csr_write                          (mm_interconnect_0_tse_0_dma_tx_prefetcher_csr_write),        //                                                     .write
		.tse_0_dma_tx_prefetcher_csr_read                           (mm_interconnect_0_tse_0_dma_tx_prefetcher_csr_read),         //                                                     .read
		.tse_0_dma_tx_prefetcher_csr_readdata                       (mm_interconnect_0_tse_0_dma_tx_prefetcher_csr_readdata),     //                                                     .readdata
		.tse_0_dma_tx_prefetcher_csr_writedata                      (mm_interconnect_0_tse_0_dma_tx_prefetcher_csr_writedata),    //                                                     .writedata
		.tse_0_tse_control_port_address                             (mm_interconnect_0_tse_0_tse_control_port_address),           //                               tse_0_tse_control_port.address
		.tse_0_tse_control_port_write                               (mm_interconnect_0_tse_0_tse_control_port_write),             //                                                     .write
		.tse_0_tse_control_port_read                                (mm_interconnect_0_tse_0_tse_control_port_read),              //                                                     .read
		.tse_0_tse_control_port_readdata                            (mm_interconnect_0_tse_0_tse_control_port_readdata),          //                                                     .readdata
		.tse_0_tse_control_port_writedata                           (mm_interconnect_0_tse_0_tse_control_port_writedata),         //                                                     .writedata
		.tse_0_tse_control_port_waitrequest                         (mm_interconnect_0_tse_0_tse_control_port_waitrequest),       //                                                     .waitrequest
		.uart_0_s1_address                                          (mm_interconnect_0_uart_0_s1_address),                        //                                            uart_0_s1.address
		.uart_0_s1_write                                            (mm_interconnect_0_uart_0_s1_write),                          //                                                     .write
		.uart_0_s1_read                                             (mm_interconnect_0_uart_0_s1_read),                           //                                                     .read
		.uart_0_s1_readdata                                         (mm_interconnect_0_uart_0_s1_readdata),                       //                                                     .readdata
		.uart_0_s1_writedata                                        (mm_interconnect_0_uart_0_s1_writedata),                      //                                                     .writedata
		.uart_0_s1_begintransfer                                    (mm_interconnect_0_uart_0_s1_begintransfer),                  //                                                     .begintransfer
		.uart_0_s1_chipselect                                       (mm_interconnect_0_uart_0_s1_chipselect)                      //                                                     .chipselect
	);

	candy_avb_test_qsys_irq_mapper irq_mapper (
		.clk           (altpll_0_c0_clk),                    //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),           // receiver6.irq
		.sender_irq    (nios2_0_irq_irq)                     //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_0_c4_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (altpll_0_c4_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	candy_avb_test_qsys_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (6),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (altpll_0_c4_clk),                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_002_reset_out_reset),    // in_rst_0.reset
		.in_0_data           (tse_0_tse_receive_data),                //     in_0.data
		.in_0_valid          (tse_0_tse_receive_valid),               //         .valid
		.in_0_ready          (tse_0_tse_receive_ready),               //         .ready
		.in_0_startofpacket  (tse_0_tse_receive_startofpacket),       //         .startofpacket
		.in_0_endofpacket    (tse_0_tse_receive_endofpacket),         //         .endofpacket
		.in_0_empty          (tse_0_tse_receive_empty),               //         .empty
		.in_0_error          (tse_0_tse_receive_error),               //         .error
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_out_0_error)          //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                    // reset_in0.reset
		.reset_in1      (nios2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                           //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_req      (),                                  // (terminated)
		.reset_req_in0  (1'b0),                              // (terminated)
		.reset_req_in1  (1'b0),                              // (terminated)
		.reset_in2      (1'b0),                              // (terminated)
		.reset_req_in2  (1'b0),                              // (terminated)
		.reset_in3      (1'b0),                              // (terminated)
		.reset_req_in3  (1'b0),                              // (terminated)
		.reset_in4      (1'b0),                              // (terminated)
		.reset_req_in4  (1'b0),                              // (terminated)
		.reset_in5      (1'b0),                              // (terminated)
		.reset_req_in5  (1'b0),                              // (terminated)
		.reset_in6      (1'b0),                              // (terminated)
		.reset_req_in6  (1'b0),                              // (terminated)
		.reset_in7      (1'b0),                              // (terminated)
		.reset_req_in7  (1'b0),                              // (terminated)
		.reset_in8      (1'b0),                              // (terminated)
		.reset_req_in8  (1'b0),                              // (terminated)
		.reset_in9      (1'b0),                              // (terminated)
		.reset_req_in9  (1'b0),                              // (terminated)
		.reset_in10     (1'b0),                              // (terminated)
		.reset_req_in10 (1'b0),                              // (terminated)
		.reset_in11     (1'b0),                              // (terminated)
		.reset_req_in11 (1'b0),                              // (terminated)
		.reset_in12     (1'b0),                              // (terminated)
		.reset_req_in12 (1'b0),                              // (terminated)
		.reset_in13     (1'b0),                              // (terminated)
		.reset_req_in13 (1'b0),                              // (terminated)
		.reset_in14     (1'b0),                              // (terminated)
		.reset_req_in14 (1'b0),                              // (terminated)
		.reset_in15     (1'b0),                              // (terminated)
		.reset_req_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_0_debug_reset_request_reset),      // reset_in1.reset
		.clk            (altpll_0_c0_clk),                        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_0_debug_reset_request_reset),  // reset_in1.reset
		.clk            (altpll_0_c4_clk),                    //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
