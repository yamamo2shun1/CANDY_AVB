��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&#;K0���r�X�	�m�q�мpN��[�#,�vJ����.	�x˰�d�������O��^�����6a�$}�.��ò�q�����\p�r�u�ۉa[%�����4%��_��Yhfʅ�gp�z8O�.�8,��]GE9;���F%C�p+�9�:�S�
)�:B��O5?�"��-f5��
��lB�^J��[�P԰w��y�� �E�Mje�]��=$s����ō5��= d��1�k;"ji0�s���h˓}���8vE9�S���5QG%Q������]�:L�-�|&H{���\����Z�zFgXMA|�P"��ð3:�R��~�`r���<��?���%�FZ��Q��7����Z�\clS���;�漩�6��q�d��SvZ�:؆Y�"%<�Fb�/ҟ�;��4|�}����Ô߿F�:w�>�J�ד�8�<m3���,�H^ߘ�be�{#O�hێ�|M�:PE�KX%��@3�䀗���u�����^4�w�j�99w:���-�P�| E����ɣ>!�w&��#&���j���l�-r>��2�������w�ʫ����@�~+< H��Y������WVȋSw�)_Z�(�r���LK���<�|�>��{�[�&�r`D��D��%Z��X4
�{�J���?ُ{k�\�W����(ԗ�劁�BXe��j9?x�9����& ځ��6x�H�D|�n��D��4�_�p��>g�d�[�̽%At3|`�;�����P�������@�qo�R���0^v�"I�J�6qI`?b��g�����%�����bdC�m����_ō%4s��a�E�����úв��2�JG�z�O���,�"<��V�MF�rCbبѣ�Q-ȱ:�5�m�D0|�#������iQ�˹�y������Y���9���UU���6�׃����o�jV��@���6�JH��3�����h�d��˅�RvC��{�oe#ՠ/
>��d�QF_��}�1�@٘Eŷ{��F������n�x��,h�(��|��xW�N@�H�Q����h���eV���PkՇ�����#�^���x^|������>?M���Z�����]K�pa���h��3�O��q��7s�ίe2R+����K�X����Г��o��u�ka?w��yəǎ�t������pN��|w"���+&,�M�ci������åEwIOr�s�+��<���LY/��*�@�w���^�ݡ�kæ�/~j�?���s<�ơ�2ܜ�U��9u_�lf4^��N���y�9(ʽx�fqk�;`�'IR�%�7)u�7�CМ�C���=D��E��H|�C1���P�9m��]�(�FDp?.�h����4}m���lF�d���%]���[�#bI S�W5!��C���ÿ�[�@g+#��IL	Yw�es[#J��(�;����:y^�a�	�&D(��R}'֟�ع`_��LX�r�Uͭ�G*(=�˙D����0k����Ł�kW_��t:ro���a�8�[���%5!����������I��]��r�K+�^)� @S?ƾM�ݵ��J#���/�XL��� � ٢�;���I��t���^V������f�Ϲ1�"d�S'Ab�0�R���j&���T���|����d�Mf��71�b����;�#�p��p���14z�l�����O�l+"�2����
�.�{�tUܐ@a�|��G6��G�� ��
CW�2�W���f0S+g���5�<����	)�WS�ZtQ�U*j�m0ʏ\-��P�T��5B�s��K���o8Y{�]�0�FL�4~B��ؽ�����'�{��ەZ�IT���5N
������j;��߽R+˼sЌT�j�h��A�9�X��*�őu�?�ic&	#�Ϊm��1t����ױ�`��Uc �H�J퐼K�6J^2jIE�����d@�����l
��N�N�����"�כ�c64�8_��>��0B�(���J&TNU��ǰ�Hl����|��@%��n�`c�լ+F�(/-G�q&I�ֶ��$�����{��:^�\L���{��^8��K9L2�����a�4Bu|?�k{��'n?H���kW���0�=D���EZ#*?Ə���&>BU|�K�%3��ʁ"�S�:�;ƸU2(X�*��;�6�[�mƱ��sk��q�r��Z��ޠ��x��w�T��gk�O�jP�<J�ۏ��tU�-�}�,�6'�j_�[@�	�a �4�@c�#%���R_��3^�!�����]�tG[����f�/�͊�'�X��PLD�	?8P"z@�0�����7M��젗���RsӖw�xӞ��#���+:��zߌ�N�8ZJ���Ti|/�>���fѮmb������-"�bF/e!��V�?�Az����3C�����%��$4m��
�K�K�\Z�a�ǡ��;K��$B��$���q��է���2j K��i�i&��vpI|��d9?�\F<�_��W[����c�ڝw\;�550{(<H�6@�"�E�!���v��ߓ�������-txZ�t����M�'{e�|���ʵ����ί����2'=��vɷ�D8 ϐ�V�����|(���Ia�Jp��k�ݿ��f9H$^��VZ���Kp!�u9%�*��r.�,=�|��-L ���?�+D�����=�xv��nk��! +�w��wCr�t(W�\��vBT�3���o��5�� ��R�
�Ydw��R͛S�a�_���R��:>�����N..��M�+�K+�]P����>���,�������-`���S?����R�æ�S<I1[h�ĉ�Z*2��A��*_G:��.���Hf'7��:�-?� �����L��`ju7��Ɨ.bg�p������;1�}�lO�#��V������Zv�*�&����D��w
]P"
��D��4���P���H��˵���v��G�e�M�p�C�g�-�#Z�?}����8͒7v>N��mRY���x@ ��?���z�^w�C� ����D3Tqa��zT}�C�(r@ZkK�����J2LPL�X����+9�����}i�>u׳����ߺ��x\���u��9�����i]�u4)�]�)���=�q��v-/j�^�Gڄ��gemg]	s|Dg����ܺr�����@�������L����e�|RBs��^C2w���~liAg�� W;D.b�$Ἆ�]m/�f�E�{�*+�Áhw�\I5EM�~�z�1��]|U��5���eB����dN�7���
!��&G��(ub� ��A@n������#��	��忀�%�ԮS��P>�2�h-qы5���� !���#� �Ђ��{LŜn�����?��Ov��lAϞ�BsL�����,�	��X����b��<���b6a��a7K3���{�{��*y�4?r� "{�Bg���߁>��1�p��������ލ�,
������� ��U9�h
ɛ�7|K�����B鉿 N��W��HE�;9u����>�+����/�VckI@�L\�*IS�O�B`�A���Ĭ���'�j�戹��K| fBN�o��l�����{�\uE�(ld4�z���*���H��pۋ
�G�@��g)��ާ�D~l�c9~�a�㔾�Ƥ��.^��'�ӱbf^31��`6v�c�oc� ��ގ�׾��P!kL������ j�#���'����z{�nߒ�����!�2u�-':I�O �����h�W�<`��@�)�Q�sv��5�2�>c��MFAu�
��.����Ya�ϯ����	�;�;�濯V�X�Ғ
0�[\�v#��i�:R(�eVs?߼]mƉaxz��3X���~�7�J� 6��n��j&��.Zc�P���\���
�{}Rf�Xj�l>OU^�tvǻ��#1�Kgĳ۽"�s/�Kk�0Θ���$cV,\����t:^�����v�عIzh�I;�-�qIX}���n�q�J9�I�~��ID5R�s�"
����! }{�RL��V�w ��>v��C֙�N���ފ������ӎ�{Ll�%=~8\�ӥ��
� �D�zƇ{҃�Bޔz�痤���p�z�Yt[f�
�� �:�/V;DՙEѸZ^�w�{`�xJ�9-#��U_H����K�	�_�Pt�	�.�8��C��-1��*�h0-�V�	쾆S�hN